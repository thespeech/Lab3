----------------------------------------------------------------------------------
-- Company: NUS
-- Engineer: Rajesh Panicker
-- 
-- Create Date:   21:06:18 14/10/2014
-- Design Name: 	PC
-- Target Devices: Nexys 4 (Artix 7 100T)
-- Tool versions: ISE 14.7
-- Description: PC for the basic MIPS processor
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: The interface (entity) as well as implementation (architecture) can be modified
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity PC is
	Port(	PC_in 	: in STD_LOGIC_VECTOR (31 downto 0);
			PC_out 	: out STD_LOGIC_VECTOR (31 downto 0) := x"00400000";
			RESET		: in STD_LOGIC;
			CLK		: in STD_LOGIC);
end PC;


architecture arch_PC of PC is
begin

--<implement PC here>

process(CLK)
begin

if (CLK'event and CLK = '1') then
	if RESET = '1' then
		PC_out <= x"00400000";
	else
		PC_out <= PC_in;
	end if;
end if;

end process;

end arch_PC;

